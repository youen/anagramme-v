module main

import vsl.iter
import os
import encoding.csv
import arrays

fn main() {
	mut anagramme := new_anagramme()
	anagramme.load_file("data/francais.txt")!
	anagramme.load_file("data/1grams_french.csv")!
	anagramme.load_file("data/2grams_french.csv")!
	anagramme.load_file("data/3grams_french.csv")!
	anagramme.load_file("data/4grams_french.csv")!
	anagramme.load_file("data/5grams_french.csv")!


//	println(anagramme.find("lino pimo")) // mini pool
//	println(anagramme.find("adrien youen")) // 'denier noyau'
//	println(anagramme.find("cgi n est pas a vendre")) // 'passant divergence'
//	println(anagramme.find("eric simon")) // roi mince
//	println(anagramme.find("france travail")) // 'flairer vacant' 
//	println(anagramme.find("cgi n est pas a vendre"))
	println(">>> ${os.args[1]}")
	for result in  anagramme.find_iterator(os.args[1]) {
		println(result)
	}
	
}

struct Anagramme {
mut:
	index map[string][]string
}

fn new_anagramme() Anagramme {
	return Anagramme{
		index : {

		}
	}
}

fn find_subseeds (seed string)  [][]string {
	ss := new_seed_splitter(seed)

	mut subseeds := [][]string{}
	for subseed in ss {
		subseeds << subseed
	}

	return subseeds

}

fn (mut a Anagramme) add( word string)  {

	a.index[a.seed(word)] << word

}

fn (mut a Anagramme) load_file(filename string) ! {
	data := os.read_file(filename) !
    mut reader := csv.new_reader(data)
	// read header
	reader.read() !
    for {
        word := reader.read() or {
            break
        }
        a.add(word[0])
    }
}

fn (a Anagramme) find( word string) []string {

	mut result :=  []string{}
	for anagramme in a.find_iterator(word) {
		result << anagramme
	}

	return arrays.distinct(result)
}

enum AnagrammeIteratorState as u8 {
	start
	direct
	subseed
	recursive
}


struct AnagrammeIterator {
	anagramme Anagramme
	seed string

mut:
	ss SeedSplitter
	state AnagrammeIteratorState
	buffer []string
	cache map[string]bool

}

fn (a Anagramme) find_iterator( word string) AnagrammeIterator {
	seed := a.seed(word)
	return AnagrammeIterator{
		anagramme : a
		seed : seed
		ss : new_seed_splitter(seed)
		state : AnagrammeIteratorState.start
	}

}

fn (mut a AnagrammeIterator) next() ?string {
	for {
		match a.state {
			.start {
				a.buffer = a.anagramme.index[a.seed]
				a.state = AnagrammeIteratorState.direct

			}
			.direct {
				if a.buffer.len > 0 {
					if a.buffer.last() in a.cache {
						a.buffer.pop()
						continue
					} else {
						result := a.buffer.pop()
						a.cache[result] = true
						return result
					}

				} else {
					a.state = AnagrammeIteratorState.subseed
				}

			}
			.subseed {
				if a.buffer.len > 0 {
		
					return a.buffer.pop()
					
				} else {
					subseed := a.ss.next() or {  
						a.state = AnagrammeIteratorState.recursive
						a.ss =  new_seed_splitter(a.seed)
						continue
					}

					first_col := a.anagramme.index[subseed[0]] or {  continue }
					second_col := a.anagramme.index[subseed[1]] or {  continue }
					for first in first_col{
						for second in second_col {
							result := "${first} ${second}"
							ratio := f64(result.count(" ")) / f64(result.len) 
							//println("${result} : ${ratio}")
							if (ratio) >  0.1 {
								continue
							}
							if !(result in a.cache ){
								a.cache[result] = true
								a.buffer <<  result
							}
						}
					}
				}

			}
			.recursive {
				if a.buffer.len > 0 {
		
					return a.buffer.pop()
					
				} else {
					subseed := a.ss.next() or { return none}

					first_col := a.anagramme.index[subseed[0]] or {  continue }
					for first in first_col{
						for second in a.anagramme.find_iterator(subseed[1]) {
							result := "${first} ${second}"
							ratio := f64(result.count(" ")) / f64(result.len) 
							if (ratio) >  0.2 {
								continue
							}
							// println("${result} : ${ratio}")
							if !(result in a.cache ){
								a.cache[result] = true
								a.buffer <<  result
							}
						}
					}
				}

			}
		}
	}
	
	return none

}

fn (a Anagramme) seed( word string) string {
	mut runes := word.replace(" ","").runes()
	runes.sort()
	return runes.string()
}

struct SeedSplitter {
	seed string
mut:
	k int
	choice_k_in ChoiceKIn
}

fn new_seed_splitter(seed string) SeedSplitter {
	return SeedSplitter {
		seed : seed,
		k : 2
		choice_k_in : new_choice_k_in(seed, 2)
	}
}

fn (mut s SeedSplitter) next() ?[]string {

	combi := s.choice_k_in.next() or { 
		if s.k < s.seed.len {
			s.k++
			s.choice_k_in = new_choice_k_in(s.seed, s.k)
			return s.next()
		}
		return none
		}

	mut first := ""
	mut second := ""
	for index in 0..s.seed.len {
		if index in combi {
			 first += s.seed[index].ascii_str()
		} else {

		second += s.seed[index].ascii_str()
		}


	}

	return [first, second]
}

struct ChoiceKIn {
mut:
	iter iter.CombinationsIter
}

fn new_choice_k_in(seed string, k int) ChoiceKIn {
	mut code := []f64{}
	for index in 0..seed.len {
		code << f64(index)
	}
	return ChoiceKIn {
		iter : iter.CombinationsIter.new(code, k)
	} 
}

fn (mut c ChoiceKIn) next() ?[]int {
	

	combi := c.iter.next() or { 
		return none
		} 

	mut combi_int := []int{}
	for n in combi {
		combi_int << int(n)
	}

	return combi_int
	
}
