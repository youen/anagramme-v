module main

fn main() {
	not_a_number := 'aa'
	number := not_a_number.int()
	println(not_a_number + number.str())	
}

fn anagramme(seed string) []string {
	return ["niche"]
}