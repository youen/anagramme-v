module main

fn test_anagrame () {
	assert "niche" in anagramme("chien")
}
